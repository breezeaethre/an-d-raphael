magic
tech sky130A
magscale 1 2
timestamp 1729416473
<< nwell >>
rect -282 -1996 516 452
rect -282 -1999 -101 -1996
rect -282 -2061 -96 -1999
rect -282 -2062 -64 -2061
rect 2 -2062 516 -1996
rect -282 -2226 516 -2062
<< nsubdiff >>
rect -246 382 -186 416
rect 420 382 480 416
rect -246 356 -212 382
rect 446 356 480 382
rect -246 -2156 -212 -2130
rect 446 -2156 480 -2130
rect -246 -2190 -186 -2156
rect 420 -2190 480 -2156
<< nsubdiffcont >>
rect -186 382 420 416
rect -246 -2130 -212 356
rect 446 -2130 480 356
rect -186 -2190 420 -2156
<< poly >>
rect -162 275 -70 291
rect -162 241 -146 275
rect -112 241 -70 275
rect -162 225 -70 241
rect -100 220 -70 225
rect 304 275 396 291
rect 304 241 346 275
rect 380 241 396 275
rect 304 225 396 241
rect 304 220 334 225
rect -162 -359 -70 -343
rect -162 -393 -146 -359
rect -112 -393 -70 -359
rect -162 -409 -70 -393
rect -100 -434 -70 -409
rect 304 -359 396 -343
rect 304 -393 346 -359
rect 380 -393 396 -359
rect 304 -409 396 -393
rect 304 -434 334 -409
rect -12 -1017 246 -757
rect -100 -1345 -70 -1340
rect -162 -1361 -70 -1345
rect -162 -1395 -146 -1361
rect -112 -1395 -70 -1361
rect -162 -1411 -70 -1395
rect 304 -1346 334 -1340
rect 304 -1362 396 -1346
rect 304 -1396 346 -1362
rect 380 -1396 396 -1362
rect 304 -1412 396 -1396
rect -100 -1999 -70 -1994
rect -162 -2015 -70 -1999
rect -162 -2049 -146 -2015
rect -112 -2049 -70 -2015
rect -162 -2065 -70 -2049
rect 304 -1999 334 -1994
rect 304 -2015 396 -1999
rect 304 -2049 346 -2015
rect 380 -2049 396 -2015
rect 304 -2065 396 -2049
<< polycont >>
rect -146 241 -112 275
rect 346 241 380 275
rect -146 -393 -112 -359
rect 346 -393 380 -359
rect -146 -1395 -112 -1361
rect 346 -1396 380 -1362
rect -146 -2049 -112 -2015
rect 346 -2049 380 -2015
<< locali >>
rect -246 382 -186 416
rect 420 382 480 416
rect -246 356 -212 382
rect 446 356 480 382
rect -162 241 -146 275
rect -112 241 -96 275
rect 330 241 346 275
rect 380 241 396 275
rect -146 181 -112 241
rect 346 179 380 241
rect -162 -393 -146 -359
rect -112 -393 -96 -359
rect 330 -393 346 -359
rect 380 -393 396 -359
rect -146 -476 -112 -393
rect -146 -1361 -112 -1302
rect -162 -1395 -146 -1361
rect -112 -1395 -96 -1361
rect 346 -1362 380 -1302
rect 330 -1396 346 -1362
rect 380 -1396 396 -1362
rect -146 -2015 -112 -1956
rect 346 -2015 380 -1956
rect -162 -2049 -146 -2015
rect -112 -2049 -96 -2015
rect 330 -2049 346 -2015
rect 380 -2049 396 -2015
rect -246 -2156 -212 -2130
rect 446 -2156 480 -2130
rect -246 -2190 -186 -2156
rect 420 -2190 480 -2156
<< viali >>
rect -146 241 -112 275
rect 346 241 380 275
rect -146 -393 -112 -359
rect 346 -393 380 -359
rect -146 -1395 -112 -1361
rect 346 -1396 380 -1362
rect -146 -2049 -112 -2015
rect 346 -2049 380 -2015
rect 88 -2190 146 -2156
<< metal1 >>
rect -158 275 -100 281
rect 334 275 392 281
rect -168 241 -146 275
rect -112 241 -82 275
rect 320 241 346 275
rect 380 241 405 275
rect -158 235 -100 241
rect 334 235 392 241
rect -184 6 -174 182
rect -122 6 -14 182
rect 79 6 89 182
rect 145 6 155 182
rect 248 6 359 182
rect 411 6 421 182
rect -6 -96 4 -44
rect 72 -96 82 -44
rect 152 -96 162 -44
rect 230 -96 240 -44
rect -158 -359 -100 -353
rect 334 -359 392 -353
rect -168 -393 -146 -359
rect -112 -393 -90 -359
rect 324 -393 346 -359
rect 380 -393 403 -359
rect -158 -399 -100 -393
rect 334 -399 392 -393
rect 345 -472 380 -399
rect -156 -648 -67 -472
rect -15 -648 -5 -472
rect 79 -648 89 -472
rect 145 -648 155 -472
rect 239 -648 249 -472
rect 301 -648 390 -472
rect 80 -741 155 -707
rect -77 -917 -71 -857
rect -11 -917 245 -857
rect 305 -917 311 -857
rect 78 -1067 155 -1033
rect -156 -1302 -67 -1126
rect -15 -1302 -5 -1126
rect 79 -1302 89 -1126
rect 145 -1302 155 -1126
rect 239 -1302 249 -1126
rect 301 -1302 390 -1126
rect -158 -1361 -100 -1355
rect -172 -1395 -146 -1361
rect -112 -1395 -92 -1361
rect 334 -1362 392 -1356
rect -158 -1401 -100 -1395
rect 324 -1396 346 -1362
rect 380 -1396 405 -1362
rect 334 -1402 392 -1396
rect -6 -1730 4 -1678
rect 72 -1730 82 -1678
rect 152 -1730 162 -1678
rect 230 -1730 240 -1678
rect -184 -1956 -174 -1780
rect -122 -1956 -14 -1780
rect 79 -1956 89 -1780
rect 145 -1956 155 -1780
rect 248 -1956 359 -1780
rect 411 -1956 422 -1780
rect -158 -2015 -100 -2009
rect 334 -2015 392 -2009
rect -168 -2049 -146 -2015
rect -112 -2049 -88 -2015
rect 320 -2049 346 -2015
rect 380 -2049 404 -2015
rect -158 -2055 -100 -2049
rect 334 -2055 392 -2049
rect 76 -2156 158 -2150
rect 76 -2190 88 -2156
rect 146 -2190 158 -2156
rect 76 -2196 158 -2190
<< via1 >>
rect -174 6 -122 182
rect 89 6 145 182
rect 359 6 411 182
rect 4 -96 72 -44
rect 162 -96 230 -44
rect -67 -648 -15 -472
rect 89 -648 145 -472
rect 249 -648 301 -472
rect -71 -917 -11 -857
rect 245 -917 305 -857
rect -67 -1302 -15 -1126
rect 89 -1302 145 -1126
rect 249 -1302 301 -1126
rect 4 -1730 72 -1678
rect 162 -1730 230 -1678
rect -174 -1956 -122 -1780
rect 89 -1956 145 -1780
rect 359 -1956 411 -1780
<< metal2 >>
rect -178 357 -118 366
rect -178 288 -118 297
rect 355 357 415 366
rect 355 288 415 297
rect -174 182 -122 288
rect -174 -1780 -122 6
rect 89 182 145 192
rect 89 -4 145 6
rect 359 182 411 288
rect -94 -35 -24 -25
rect 4 -42 230 -34
rect 4 -44 266 -42
rect -24 -96 4 -44
rect 72 -96 162 -44
rect 230 -96 266 -44
rect -94 -115 -24 -105
rect 4 -98 266 -96
rect 322 -98 331 -42
rect 4 -106 230 -98
rect -67 -472 -15 -462
rect 89 -472 145 -462
rect 249 -472 301 -462
rect -77 -857 -5 -648
rect 89 -658 145 -648
rect -77 -917 -71 -857
rect -11 -917 -5 -857
rect -77 -1126 -5 -917
rect 239 -857 311 -648
rect 239 -917 245 -857
rect 305 -917 311 -857
rect 89 -1126 145 -1116
rect 239 -1126 311 -917
rect -67 -1312 -15 -1302
rect 89 -1312 145 -1302
rect 249 -1312 301 -1302
rect -87 -1674 -31 -1667
rect 4 -1674 230 -1668
rect -89 -1676 230 -1674
rect -89 -1732 -87 -1676
rect -31 -1678 230 -1676
rect 259 -1669 329 -1659
rect -31 -1730 4 -1678
rect 72 -1730 162 -1678
rect 230 -1730 259 -1678
rect -31 -1732 230 -1730
rect -89 -1734 230 -1732
rect -87 -1741 -31 -1734
rect 4 -1740 230 -1734
rect 259 -1749 329 -1739
rect -174 -2062 -122 -1956
rect 89 -1780 145 -1770
rect 89 -1966 145 -1956
rect 359 -1780 411 6
rect 359 -2062 411 -1956
rect -178 -2071 -118 -2062
rect -178 -2140 -118 -2131
rect 355 -2071 415 -2062
rect 355 -2140 415 -2131
<< via2 >>
rect -178 297 -118 357
rect 355 297 415 357
rect 89 6 145 182
rect -94 -105 -24 -35
rect 266 -98 322 -42
rect 89 -648 145 -472
rect 89 -1302 145 -1126
rect -87 -1732 -31 -1676
rect 259 -1739 329 -1669
rect 89 -1956 145 -1780
rect -178 -2131 -118 -2071
rect 355 -2131 415 -2071
<< metal3 >>
rect -183 357 -113 362
rect 350 357 420 362
rect -183 297 -178 357
rect -118 297 355 357
rect 415 297 420 357
rect -183 292 -113 297
rect 350 292 420 297
rect 79 182 155 187
rect 79 6 89 182
rect 145 6 155 182
rect -104 -35 -14 -30
rect -104 -105 -94 -35
rect -24 -105 -14 -35
rect -104 -110 -14 -105
rect -89 -1671 -29 -110
rect 79 -472 155 6
rect 261 -42 327 -37
rect 261 -98 266 -42
rect 322 -98 327 -42
rect 261 -103 327 -98
rect 79 -648 89 -472
rect 145 -648 155 -472
rect 79 -1126 155 -648
rect 79 -1302 89 -1126
rect 145 -1302 155 -1126
rect -92 -1676 -26 -1671
rect -92 -1732 -87 -1676
rect -31 -1732 -26 -1676
rect -92 -1737 -26 -1732
rect 79 -1780 155 -1302
rect 264 -1664 324 -103
rect 249 -1669 339 -1664
rect 249 -1739 259 -1669
rect 329 -1739 339 -1669
rect 249 -1744 339 -1739
rect 79 -1956 89 -1780
rect 145 -1956 155 -1780
rect 79 -1961 155 -1956
rect -183 -2071 -113 -2066
rect 350 -2071 420 -2066
rect -183 -2131 -178 -2071
rect -118 -2131 355 -2071
rect 415 -2131 420 -2071
rect -183 -2136 -113 -2131
rect 350 -2136 420 -2131
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729416473
transform 1 0 -85 0 1 -560
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729416473
transform 1 0 -85 0 1 -1868
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729416473
transform 1 0 -85 0 1 94
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729416473
transform 1 0 319 0 1 94
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729416473
transform 1 0 319 0 1 -560
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729416473
transform 1 0 319 0 1 -1214
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729416473
transform 1 0 -85 0 1 -1214
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729416473
transform 1 0 319 0 1 -1868
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_0
timestamp 1729396642
transform 1 0 117 0 1 -1868
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_1
timestamp 1729396642
transform 1 0 117 0 1 94
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_2
timestamp 1729396642
transform 1 0 117 0 1 -560
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_3
timestamp 1729396642
transform 1 0 117 0 1 -1214
box -223 -200 223 200
<< labels >>
flabel nwell 36 -1868 36 -1868 0 FreeSans 160 0 0 0 M7
flabel nwell 200 -1867 200 -1867 0 FreeSans 160 0 0 0 M7
flabel nwell 34 -1215 34 -1215 0 FreeSans 160 0 0 0 M6
flabel nwell 201 -1212 201 -1212 0 FreeSans 160 0 0 0 M6
flabel nwell 33 -560 33 -560 0 FreeSans 160 0 0 0 M6
flabel nwell 196 -560 196 -560 0 FreeSans 160 0 0 0 M6
flabel metal1 83 -2172 83 -2172 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal3 114 -1525 114 -1525 0 FreeSans 800 0 0 0 D5
port 2 nsew
flabel metal1 115 -1051 115 -1051 0 FreeSans 800 0 0 0 VIN
port 3 nsew
flabel metal1 323 -1210 323 -1210 0 FreeSans 800 0 0 0 D6
port 4 nsew
flabel metal2 112 -69 112 -69 0 FreeSans 800 0 0 0 VIP
port 6 nsew
flabel metal1 -87 99 -87 99 0 FreeSans 800 0 0 0 OUT
port 5 nsew
flabel nwell 201 92 201 92 0 FreeSans 160 0 0 0 M7
flabel nwell 34 95 34 95 0 FreeSans 160 0 0 0 M7
<< end >>
