magic
tech sky130A
magscale 1 2
timestamp 1729430370
<< viali >>
rect -60 3362 -26 3396
rect -473 1374 -425 1408
<< metal1 >>
rect -72 3396 56 3408
rect -72 3362 -60 3396
rect -26 3362 56 3396
rect -72 3350 56 3362
rect 820 2184 1069 2230
rect -1509 2016 -788 2050
rect -1509 -36 -1475 2016
rect -791 1534 -781 1586
rect -729 1534 -719 1586
rect -87 1479 182 1525
rect -473 1414 -426 1462
rect -485 1408 -413 1414
rect -485 1374 -473 1408
rect -425 1374 -413 1408
rect -485 1368 -413 1374
rect -1358 693 -1348 745
rect -1296 741 -1286 745
rect -1296 696 -690 741
rect -1296 693 -1286 696
rect -87 657 -41 1479
rect 17 793 23 845
rect 75 793 184 845
rect -412 611 -41 657
rect 741 17 817 139
rect -1509 -70 -813 -36
rect -847 -170 -813 -70
rect 278 -59 817 17
rect 278 -361 354 -59
rect 268 -437 278 -361
rect 354 -437 364 -361
rect -199 -878 -153 -511
<< via1 >>
rect -781 1534 -729 1586
rect -1348 693 -1296 745
rect 23 793 75 845
rect 278 -437 354 -361
<< metal2 >>
rect -781 1586 -729 1596
rect -1517 1534 -781 1586
rect -1517 -159 -1465 1534
rect -781 1524 -729 1534
rect 23 845 75 851
rect -1352 749 -1292 759
rect 23 745 75 793
rect -415 693 75 745
rect -1352 679 -1292 689
rect 278 -361 354 -351
rect 278 -447 354 -437
rect -1063 -877 -1011 -641
<< via2 >>
rect -1352 745 -1292 749
rect -1352 693 -1348 745
rect -1348 693 -1296 745
rect -1296 693 -1292 745
rect -1352 689 -1292 693
rect 278 -437 354 -361
<< metal3 >>
rect -1362 749 -1282 754
rect -1641 689 -1352 749
rect -1292 689 -1282 749
rect -1362 684 -1282 689
rect 268 -361 364 -356
rect 268 -437 278 -361
rect 354 -437 364 -361
rect 268 -442 364 -437
rect 287 -868 347 -546
use nmoscs34  nmoscs34_0
timestamp 1729333487
transform 1 0 -656 0 1 765
box -770 -745 630 649
use nmoscs89  nmoscs89_0
timestamp 1729423161
transform 1 0 -696 0 1 2952
box -176 -1496 670 445
use pmoscs67  pmoscs67_0
timestamp 1729416473
transform 0 1 548 -1 0 -282
box -282 -2226 516 452
use pmoscs  pmoscs_0
timestamp 1729237752
transform 1 0 153 0 1 1705
box -153 -1705 846 1155
<< labels >>
flabel metal1 1042 2210 1042 2210 0 FreeSans 480 0 0 0 VDD_OA
port 0 nsew
flabel metal1 21 3382 21 3382 0 FreeSans 480 0 0 0 GND_OA
port 1 nsew
flabel metal3 -1587 721 -1587 721 0 FreeSans 480 0 0 0 RS_OA
port 2 nsew
flabel metal1 -180 -845 -180 -845 0 FreeSans 480 0 0 0 VIN_OA
port 3 nsew
flabel metal3 319 -837 319 -837 0 FreeSans 480 0 0 0 VIP_OA
port 4 nsew
flabel metal2 -1044 -846 -1044 -846 0 FreeSans 480 0 0 0 OUT_OA
port 5 nsew
<< end >>
