** sch_path: /home/raphael03/MSIB/Inverter/ring_osc.sch
**.subckt ring_osc vdd out gnd
*.opin out
*.iopin vdd
*.iopin gnd
x1 vdd net1 out gnd inverter
x2 vdd net2 net1 gnd inverter
x3 vdd out net2 gnd inverter
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/raphael03/MSIB/Inverter/inverter.sym
** sch_path: /home/raphael03/MSIB/Inverter/inverter.sch

.end
