magic
tech sky130A
magscale 1 2
timestamp 1729237752
<< nwell >>
rect -153 -1705 846 1155
<< nsubdiff >>
rect -117 1085 -57 1119
rect 750 1085 810 1119
rect -117 1059 -83 1085
rect 776 1059 810 1085
rect -117 -1635 -83 -1609
rect 776 -1635 810 -1609
rect -117 -1669 -57 -1635
rect 750 -1669 810 -1635
<< nsubdiffcont >>
rect -57 1085 750 1119
rect -117 -1609 -83 1059
rect 776 -1609 810 1059
rect -57 -1669 750 -1635
<< poly >>
rect -33 1047 59 1063
rect -33 1013 -17 1047
rect 17 1013 59 1047
rect -33 997 59 1013
rect 29 966 59 997
rect 633 1047 725 1063
rect 633 1013 675 1047
rect 709 1013 725 1047
rect 633 997 725 1013
rect 633 991 663 997
rect 117 369 318 470
rect 634 353 726 369
rect 634 319 676 353
rect 710 319 726 353
rect 634 303 726 319
rect 634 272 664 303
rect 30 -159 60 -128
rect -32 -175 60 -159
rect -32 -209 -16 -175
rect 18 -209 60 -175
rect -32 -225 60 -209
rect 118 -325 576 -225
rect 30 -853 60 -822
rect -32 -869 60 -853
rect -32 -903 -16 -869
rect 18 -903 60 -869
rect -32 -919 60 -903
rect 634 -853 664 -822
rect 634 -869 726 -853
rect 634 -903 676 -869
rect 710 -903 726 -869
rect 376 -1021 576 -918
rect 634 -919 726 -903
rect 30 -1547 60 -1516
rect -32 -1563 60 -1547
rect -32 -1597 -16 -1563
rect 18 -1597 60 -1563
rect -32 -1613 60 -1597
rect 634 -1547 664 -1516
rect 634 -1563 726 -1547
rect 634 -1597 676 -1563
rect 710 -1597 726 -1563
rect 634 -1613 726 -1597
<< polycont >>
rect -17 1013 17 1047
rect 675 1013 709 1047
rect 676 319 710 353
rect -16 -209 18 -175
rect -16 -903 18 -869
rect 676 -903 710 -869
rect -16 -1597 18 -1563
rect 676 -1597 710 -1563
<< locali >>
rect -117 1085 -57 1119
rect 750 1085 810 1119
rect -117 1059 -83 1085
rect 776 1059 810 1085
rect -33 1013 -17 1047
rect 17 1013 33 1047
rect 659 1013 675 1047
rect 709 1013 725 1047
rect -17 966 17 1013
rect 71 966 105 970
rect 675 954 709 1013
rect 660 319 676 353
rect 710 319 726 353
rect 588 272 622 276
rect 676 272 710 319
rect -16 -175 18 -128
rect 72 -132 106 -128
rect -32 -209 -16 -175
rect 18 -209 34 -175
rect -16 -869 18 -822
rect 72 -826 106 -822
rect 588 -826 622 -822
rect 676 -869 710 -822
rect -32 -903 -16 -869
rect 18 -903 34 -869
rect 660 -903 676 -869
rect 710 -903 726 -869
rect -16 -1563 18 -1516
rect 72 -1520 106 -1516
rect 588 -1520 622 -1516
rect 676 -1563 710 -1516
rect -32 -1597 -16 -1563
rect 18 -1597 34 -1563
rect 660 -1597 676 -1563
rect 710 -1597 726 -1563
rect -117 -1635 -83 -1609
rect 776 -1635 810 -1609
rect -117 -1669 -57 -1635
rect 750 -1669 810 -1635
<< viali >>
rect -17 1013 17 1047
rect 675 1013 709 1047
rect 776 1012 810 1046
rect 676 319 710 353
rect -16 -209 18 -175
rect -16 -903 18 -869
rect 676 -903 710 -869
rect -16 -1597 18 -1563
rect 676 -1597 710 -1563
<< metal1 >>
rect -29 1047 29 1053
rect 663 1052 721 1053
rect 663 1047 823 1052
rect -29 1013 -17 1047
rect 17 1013 105 1047
rect -29 1007 29 1013
rect -17 966 17 1007
rect 71 966 105 1013
rect 587 1013 675 1047
rect 709 1046 823 1047
rect 709 1013 776 1046
rect -36 578 -26 954
rect 26 578 36 954
rect 324 525 369 966
rect 587 961 621 1013
rect 663 1012 776 1013
rect 810 1012 823 1046
rect 663 1007 823 1012
rect 664 1006 823 1007
rect 675 954 709 1006
rect 581 525 627 566
rect 669 525 715 566
rect 324 479 404 525
rect 546 479 715 525
rect -16 -169 18 -128
rect -28 -175 30 -169
rect 66 -175 112 -128
rect -28 -209 -16 -175
rect 18 -209 112 -175
rect -28 -215 30 -209
rect 66 -250 112 -209
rect 53 -302 63 -250
rect 115 -302 125 -250
rect 66 -381 147 -335
rect 66 -422 113 -381
rect -22 -822 112 -422
rect -16 -863 18 -822
rect -28 -869 30 -863
rect 72 -869 106 -822
rect -28 -903 -16 -869
rect 18 -903 106 -869
rect -28 -909 30 -903
rect 324 -1029 369 479
rect 664 353 722 359
rect 588 319 676 353
rect 710 319 722 353
rect 588 272 622 319
rect 664 313 722 319
rect 676 272 710 313
rect 582 -128 716 272
rect 582 -169 628 -128
rect 547 -215 628 -169
rect 573 -302 579 -250
rect 631 -302 637 -250
rect 582 -429 628 -302
rect 588 -869 622 -822
rect 676 -863 710 -822
rect 664 -869 722 -863
rect 588 -903 676 -869
rect 710 -903 722 -869
rect 664 -909 722 -903
rect -22 -1075 147 -1029
rect 289 -1075 369 -1029
rect -22 -1116 24 -1075
rect 66 -1116 112 -1075
rect 324 -1516 369 -1075
rect 657 -1504 667 -1128
rect 719 -1504 729 -1128
rect -16 -1557 18 -1516
rect -28 -1563 30 -1557
rect 72 -1563 106 -1516
rect -28 -1597 -16 -1563
rect 18 -1597 106 -1563
rect 588 -1563 622 -1516
rect 676 -1557 710 -1516
rect 664 -1563 722 -1557
rect 588 -1597 676 -1563
rect 710 -1597 722 -1563
rect -28 -1603 30 -1597
rect 664 -1603 722 -1597
<< via1 >>
rect -26 578 26 954
rect 63 -302 115 -250
rect 579 -302 631 -250
rect 667 -1504 719 -1128
<< metal2 >>
rect -26 954 26 964
rect -30 578 -26 625
rect 26 578 30 625
rect -30 453 30 578
rect -30 449 31 453
rect -30 393 -28 449
rect 28 393 31 449
rect -30 391 31 393
rect 654 391 663 451
rect 723 391 732 451
rect -29 -941 31 391
rect 63 -250 115 -240
rect 579 -250 631 -244
rect 115 -299 579 -253
rect 63 -312 115 -302
rect 579 -308 631 -302
rect 667 -939 719 391
rect -36 -997 -27 -941
rect 29 -997 38 -941
rect -29 -999 31 -997
rect 654 -999 663 -939
rect 723 -999 732 -939
rect 667 -1128 719 -999
rect 667 -1514 719 -1504
<< via2 >>
rect -28 393 28 449
rect 663 391 723 451
rect -27 -997 29 -941
rect 663 -999 723 -939
<< metal3 >>
rect -33 451 33 454
rect 658 451 728 456
rect -33 449 663 451
rect -33 393 -28 449
rect 28 393 663 449
rect -33 391 663 393
rect 723 391 728 451
rect -33 388 33 391
rect 658 386 728 391
rect -32 -939 34 -936
rect 658 -939 728 -934
rect -32 -941 663 -939
rect -32 -997 -27 -941
rect 29 -997 663 -941
rect -32 -999 663 -997
rect 723 -999 728 -939
rect -32 -1002 34 -999
rect 658 -1004 728 -999
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729133638
transform 1 0 45 0 1 -1316
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729133638
transform 1 0 45 0 1 -622
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729133638
transform 1 0 45 0 1 72
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729133638
transform 1 0 44 0 1 766
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729133638
transform 1 0 649 0 1 -1316
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729133638
transform 1 0 648 0 1 766
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729133638
transform 1 0 649 0 1 72
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_8
timestamp 1729133638
transform 1 0 649 0 1 -622
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729143223
transform 1 0 346 0 1 766
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729143223
transform 1 0 347 0 1 72
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729143223
transform 1 0 347 0 1 -622
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729143223
transform 1 0 347 0 1 -1316
box -323 -300 323 300
<< labels >>
flabel metal1 594 -378 594 -378 0 FreeSans 800 0 0 0 D1
port 0 nsew
flabel metal1 598 -1536 598 -1536 0 FreeSans 800 0 0 0 D5
port 1 nsew
flabel metal1 606 290 606 290 0 FreeSans 800 0 0 0 D2
port 2 nsew
flabel metal1 594 1022 594 1022 0 FreeSans 800 0 0 0 VDD
port 3 nsew
<< end >>
