magic
tech sky130A
magscale 1 2
timestamp 1728979425
<< error_p >>
rect -29 -107 29 -101
rect -29 -141 -17 -107
rect -29 -147 29 -141
<< pwell >>
rect -211 -279 211 279
<< nmos >>
rect -15 -69 15 131
<< ndiff >>
rect -73 119 -15 131
rect -73 -57 -61 119
rect -27 -57 -15 119
rect -73 -69 -15 -57
rect 15 119 73 131
rect 15 -57 27 119
rect 61 -57 73 119
rect 15 -69 73 -57
<< ndiffc >>
rect -61 -57 -27 119
rect 27 -57 61 119
<< psubdiff >>
rect -175 209 -79 243
rect 79 209 175 243
rect -175 147 -141 209
rect 141 147 175 209
rect -175 -209 -141 -147
rect 141 -209 175 -147
rect -175 -243 -79 -209
rect 79 -243 175 -209
<< psubdiffcont >>
rect -79 209 79 243
rect -175 -147 -141 147
rect 141 -147 175 147
rect -79 -243 79 -209
<< poly >>
rect -15 131 15 157
rect -15 -91 15 -69
rect -33 -107 33 -91
rect -33 -141 -17 -107
rect 17 -141 33 -107
rect -33 -157 33 -141
<< polycont >>
rect -17 -141 17 -107
<< locali >>
rect -175 209 -79 243
rect 79 209 175 243
rect -175 147 -141 209
rect 141 147 175 209
rect -61 119 -27 135
rect -61 -73 -27 -57
rect 27 119 61 135
rect 27 -73 61 -57
rect -33 -141 -17 -107
rect 17 -141 33 -107
rect -175 -209 -141 -147
rect 141 -209 175 -147
rect -175 -243 -79 -209
rect 79 -243 175 -209
<< viali >>
rect -61 -57 -27 119
rect 27 -57 61 119
rect -17 -141 17 -107
<< metal1 >>
rect -67 119 -21 131
rect -67 -57 -61 119
rect -27 -57 -21 119
rect -67 -69 -21 -57
rect 21 119 67 131
rect 21 -57 27 119
rect 61 -57 67 119
rect 21 -69 67 -57
rect -29 -107 29 -101
rect -29 -141 -17 -107
rect 17 -141 29 -107
rect -29 -147 29 -141
<< properties >>
string FIXED_BBOX -158 -226 158 226
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
