magic
tech sky130A
magscale 1 2
timestamp 1729404826
<< error_p >>
rect -108 181 -50 187
rect 50 181 108 187
rect -108 147 -96 181
rect 50 147 62 181
rect -108 141 -50 147
rect 50 141 108 147
rect -108 -147 -50 -141
rect 50 -147 108 -141
rect -108 -181 -96 -147
rect 50 -181 62 -147
rect -108 -187 -50 -181
rect 50 -187 108 -181
<< nwell >>
rect -223 -200 223 200
<< pmos >>
rect -129 -100 -29 100
rect 29 -100 129 100
<< pdiff >>
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
<< pdiffc >>
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
<< poly >>
rect -129 181 -29 197
rect -129 147 -113 181
rect -45 147 -29 181
rect -129 100 -29 147
rect 29 181 129 197
rect 29 147 45 181
rect 113 147 129 181
rect 29 100 129 147
rect -129 -147 -29 -100
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect -129 -197 -29 -181
rect 29 -147 129 -100
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 29 -197 129 -181
<< polycont >>
rect -113 147 -45 181
rect 45 147 113 181
rect -113 -181 -45 -147
rect 45 -181 113 -147
<< locali >>
rect -129 147 -113 181
rect -45 147 -29 181
rect 29 147 45 181
rect 113 147 129 181
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 113 -181 129 -147
<< viali >>
rect -96 147 -62 181
rect 62 147 96 181
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect -96 -181 -62 -147
rect 62 -181 96 -147
<< metal1 >>
rect -108 181 -50 187
rect -108 147 -96 181
rect -62 147 -50 181
rect -108 141 -50 147
rect 50 181 108 187
rect 50 147 62 181
rect 96 147 108 181
rect 50 141 108 147
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect -108 -147 -50 -141
rect -108 -181 -96 -147
rect -62 -181 -50 -147
rect -108 -187 -50 -181
rect 50 -147 108 -141
rect 50 -181 62 -147
rect 96 -181 108 -147
rect 50 -187 108 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 30 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
