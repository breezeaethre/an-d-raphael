magic
tech sky130A
magscale 1 2
timestamp 1729245583
<< nwell >>
rect -438 -1241 -122 1241
<< pwell >>
rect -705 1241 705 1507
rect -705 -1241 -438 1241
rect -122 -1241 705 1241
rect -705 -1507 705 -1241
<< mvnmos >>
rect 37 109 249 1109
rect 37 -1109 249 -109
<< mvndiff >>
rect 249 1097 307 1109
rect 249 121 261 1097
rect 295 121 307 1097
rect 249 109 307 121
rect 249 -121 307 -109
rect 249 -1097 261 -121
rect 295 -1097 307 -121
rect 249 -1109 307 -1097
<< mvndiffc >>
rect 261 121 295 1097
rect 261 -1097 295 -121
<< mvpsubdiff >>
rect -669 1459 669 1471
rect -669 1425 -561 1459
rect 561 1425 669 1459
rect -669 1413 669 1425
rect -669 1363 -611 1413
rect -669 -1363 -657 1363
rect -623 -1363 -611 1363
rect 611 1363 669 1413
rect -669 -1413 -611 -1363
rect 611 -1363 623 1363
rect 657 -1363 669 1363
rect 611 -1413 669 -1363
rect -669 -1425 669 -1413
rect -669 -1459 -561 -1425
rect 561 -1459 669 -1425
rect -669 -1471 669 -1459
<< mvnsubdiff >>
rect -306 1085 -254 1109
rect -306 133 -297 1085
rect -263 133 -254 1085
rect -306 109 -254 133
rect -306 -133 -254 -109
rect -306 -1085 -297 -133
rect -263 -1085 -254 -133
rect -306 -1109 -254 -1085
<< mvpsubdiffcont >>
rect -561 1425 561 1459
rect -657 -1363 -623 1363
rect 623 -1363 657 1363
rect -561 -1459 561 -1425
<< mvnsubdiffcont >>
rect -297 133 -263 1085
rect -297 -1085 -263 -133
<< extdrain >>
rect -254 109 37 1109
rect -254 -1109 37 -109
<< poly >>
rect 37 1181 249 1197
rect 37 1147 53 1181
rect 233 1147 249 1181
rect 37 1109 249 1147
rect 37 71 249 109
rect 37 37 53 71
rect 233 37 249 71
rect 37 21 249 37
rect 37 -37 249 -21
rect 37 -71 53 -37
rect 233 -71 249 -37
rect 37 -109 249 -71
rect 37 -1147 249 -1109
rect 37 -1181 53 -1147
rect 233 -1181 249 -1147
rect 37 -1197 249 -1181
<< polycont >>
rect 53 1147 233 1181
rect 53 37 233 71
rect 53 -71 233 -37
rect 53 -1181 233 -1147
<< locali >>
rect -657 1425 -561 1459
rect 561 1425 657 1459
rect -657 1363 -623 1425
rect 623 1363 657 1425
rect 37 1147 53 1181
rect 233 1147 249 1181
rect -297 1097 -263 1101
rect -297 117 -263 121
rect 261 1097 295 1113
rect 261 105 295 121
rect 37 37 53 71
rect 233 37 249 71
rect 37 -71 53 -37
rect 233 -71 249 -37
rect -297 -121 -263 -117
rect -297 -1101 -263 -1097
rect 261 -121 295 -105
rect 261 -1113 295 -1097
rect 37 -1181 53 -1147
rect 233 -1181 249 -1147
rect -657 -1425 -623 -1363
rect 623 -1425 657 -1363
rect -657 -1459 -561 -1425
rect 561 -1459 657 -1425
<< viali >>
rect 53 1147 233 1181
rect -297 1085 -263 1097
rect -297 133 -263 1085
rect -297 121 -263 133
rect 261 121 295 1097
rect 53 37 233 71
rect 53 -71 233 -37
rect -297 -133 -263 -121
rect -297 -1085 -263 -133
rect -297 -1097 -263 -1085
rect 261 -1097 295 -121
rect 53 -1181 233 -1147
<< metal1 >>
rect 41 1181 245 1187
rect 41 1147 53 1181
rect 233 1147 245 1181
rect 41 1141 245 1147
rect -303 1097 -257 1109
rect -303 121 -297 1097
rect -263 121 -257 1097
rect -303 109 -257 121
rect 255 1097 301 1109
rect 255 121 261 1097
rect 295 121 301 1097
rect 255 109 301 121
rect 41 71 245 77
rect 41 37 53 71
rect 233 37 245 71
rect 41 31 245 37
rect 41 -37 245 -31
rect 41 -71 53 -37
rect 233 -71 245 -37
rect 41 -77 245 -71
rect -303 -121 -257 -109
rect -303 -1097 -297 -121
rect -263 -1097 -257 -121
rect -303 -1109 -257 -1097
rect 255 -121 301 -109
rect 255 -1097 261 -121
rect 295 -1097 301 -121
rect 255 -1109 301 -1097
rect 41 -1147 245 -1141
rect 41 -1181 53 -1147
rect 233 -1181 245 -1147
rect 41 -1187 245 -1181
<< properties >>
string FIXED_BBOX -640 -1442 640 1442
string gencell sky130_fd_pr__nfet_g5v0d16v0
string library sky130
string parameters w 5.00 l 1.055 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 1.050 wmin 5.00 full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
